library verilog;
use verilog.vl_types.all;
entity FancyRegister_vlg_check_tst is
    port(
        q0              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FancyRegister_vlg_check_tst;
