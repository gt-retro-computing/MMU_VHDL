library verilog;
use verilog.vl_types.all;
entity FancyRegister_vlg_vec_tst is
end FancyRegister_vlg_vec_tst;
